interface intf();
  
  logic rst;
  logic clk;
  logic count;
  logic out;
  
endinterface
