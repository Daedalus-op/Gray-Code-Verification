`include "transaction.sv"
`include "generator.sv"
`include "driver.sv"
`include "monitor.sv"
`include "scoreboard.sv"

class environment;
	generator 	gen;
	driver    	driv;
	monitor   	mon;
	scoreboard	scb;
	mailbox 		m1;
	mailbox 		m2;

	virtual intf vif;
	function new(virtual intf vif);
		this.vif = vif;
		m1   = new();
		m2   = new();
		gen  = new(m1);
		driv = new(vif,m1);
		mon  = new(vif,m2);
		scb  = new(m2);
	endfunction
	
	task gener();
		fork 
			$display("xxxxxxxx Generating xxxxxxxx");
			gen.main();
		join
	endtask
	
	task test();
		fork
			$display("xxxxxxxxxx Testing xxxxxxxxxx");
			driv.main();
			mon.main();
			scb.main();
		join
	endtask

	
	task run;
		gener();
		repeat(4) begin
			#1;
			test();
		end
		$finish;
	endtask
	
endclass
