interface intf();

	logic rst;
	logic clk;
	logic [3:0] count;
	logic [3:0] out;

endinterface
